module pac_ROM(
    clk,
    x,
    y,
    direction,
    pixel
);

input clk;
input [4:0] x,y;
input [3:0] direction;

output reg pixel;

reg [23: 0] counter;
reg flag;


localparam L = 4'b1000;
localparam U = 4'b0100;
localparam R = 4'b0010;
localparam D = 4'b0001;



    localparam PAC_RIGHT = {
        16'b0000011111100000,
        16'b0000111111110000,
        16'b0001111111111100,
        16'b0011111111111100,
        16'b0011111111111110,
        16'b0000111111111110,
        16'b0000000111111111,
        16'b0000000000111111,
        16'b0000000000111111,
        16'b0000000111111111,
        16'b0000111111111110,
        16'b0011111111111110,
        16'b0011111111111100,
        16'b0001111111111100,
        16'b0000111111110000,
        16'b0000001111000000
        };

        localparam PAC_RIGHT_WIDE = {
            16'b0000011111100000,
            16'b0000111111110000,
            16'b0000011111111100,
            16'b0000001111111100,
            16'b0000000111111110,
            16'b0000000011111110,
            16'b0000000001111111,
            16'b0000000000111111,
            16'b0000000000111111,
            16'b0000000001111111,
            16'b0000000011111110,
            16'b0000000111111110,
            16'b0000001111111100,
            16'b0000011111111100,
            16'b0000111111110000,
            16'b0000001111000000
        };

    localparam PAC_LEFT = {
        16'b0000011111100000,
        16'b0000111111110000,
        16'b0011111111111000,
        16'b0011111111111100,
        16'b0111111111111100,
        16'b1111111111110000,
        16'b1111111110000000,
        16'b1111110000000000,
        16'b1111110000000000,
        16'b1111111110000000,
        16'b1111111111110000,
        16'b0111111111111100,
        16'b0011111111111100,
        16'b0011111111111000,
        16'b0000111111110000,
        16'b0000001111000000
        };

        localparam PAC_LEFT_WIDE = {
            16'b0000011111100000,
            16'b0000111111110000,
            16'b0011111111100000,
            16'b0011111111000000,
            16'b0111111110000000,
            16'b1111111100000000,
            16'b1111111000000000,
            16'b1111110000000000,
            16'b1111110000000000,
            16'b1111111000000000,
            16'b1111111100000000,
            16'b0111111110000000,
            16'b0011111111000000,
            16'b0011111111100000,
            16'b0000111111110000,
            16'b0000001111000000
            };

            localparam PAC_UP = {
                16'b0000000000000000,
                16'b0000000000000000,
                16'b0001100000011000,
                16'b0011100000011100,
                16'b0111110000111110,
                16'b1111110000111110,
                16'b1111110000111111,
                16'b1111111001111111,
                16'b1111111001111111,
                16'b1111111001111111,
                16'b1111111111111110,
                16'b0111111111111110,
                16'b0011111111111100,
                16'b0011111111111100,
                16'b0000111111110000,
                16'b0000001111000000
                };

            localparam PAC_UP_WIDE = {

                16'b0000000000000000,
                16'b0000000000000000,
                16'b0000000000000000,
                16'b0000000000000000,
                16'b0000000000000000,
                16'b0110000000000110,
                16'b1111000000001111,
                16'b1111100000011111,
                16'b1111110000111111,
                16'b1111111001111111,
                16'b1111111111111110,
                16'b0111111111111110,
                16'b0011111111111100,
                16'b0011111111111100,
                16'b0000111111110000,
                16'b0000001111000000
                };

            localparam PAC_DOWN = {

                16'b0000011111100000,
                16'b0000111111110000,
                16'b0011111111111100,
                16'b0011111111111100,
                16'b0111111111111110,
                16'b1111111111111110,
                16'b1111111001111111,
                16'b1111111001111111,
                16'b1111111001111111,
                16'b1111110000111111,
                16'b1111110000111110,
                16'b0111110000111110,
                16'b0011100000011100,
                16'b0001100000011000,
                16'b0000000000000000,
                16'b0000000000000000
                };

                localparam PAC_DOWN_WIDE = {

                    16'b0000011111100000,
                    16'b0000111111110000,
                    16'b0011111111111100,
                    16'b0011111111111100,
                    16'b0111111111111110,
                    16'b1111111111111110,
                    16'b1111111001111111,
                    16'b1111110000111111,
                    16'b1111100000011111,
                    16'b1111000000001111,
                    16'b0110000000000110,
                    16'b0000000000000000,
                    16'b0000000000000000,
                    16'b0000000000000000,
                    16'b0000000000000000,
                    16'b0000000000000000
                    };


    initial begin
        counter = 0;
        flag = 0;
    end

    always @(posedge clk)
    begin
        if (counter == 10000000)
        begin
            counter <= 0;
            flag <= ~flag;
        end
        else
            counter <= counter + 1;
    end

    always @(posedge clk)
    begin
        case (direction)
            L:
            begin
                if (flag)
                    pixel <= PAC_LEFT[(y / 3) * 2 * 12 + (x / 3) * 2];
                else
                    pixel <= PAC_LEFT_WIDE[(y/3) * 2 * 12 + (x/ 3) * 2];
            end
            U:
            begin
                if (flag)
                    pixel <= PAC_UP[(y / 3) * 2 * 12 + (x / 3) * 2];
                else
                    pixel <= PAC_UP_WIDE[(y/3) * 2 * 12 + (x/3) * 2];
            end
            R:
            begin
                if (flag)
                    pixel <= PAC_RIGHT[(y / 3) * 2 * 12 + (x / 3) * 2];
                else
                    pixel <= PAC_RIGHT_WIDE[(y / 3) * 2 * 12 + (x / 3) * 2];
            end
            D:
            begin
                if (flag)
                    pixel <= PAC_DOWN[(y / 3) * 2 * 12 + (x / 3) * 2];
                else
                    pixel <= PAC_DOWN_WIDE[(y / 3) * 2 * 12 + ( x / 3) * 2];
            end
            default: 
            begin
                pixel <= PAC_RIGHT[(y/3) * 2 * 12 + (x/3) * 2];
            end
        endcase
    end

endmodule

