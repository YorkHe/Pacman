`timescale 1ns/1ps

module dotMap(
    clk,
    set_x,
    set_y,
    query_x,
    query_y,
    dot,
    new
);

input clk;
input [10:0] set_x, set_y, query_x, query_y;

output dot;
output reg new;

reg[1:0] map[29*34:0];

initial begin
    map[0]=0;
    map[1]=0;
    map[2]=0;
    map[3]=0;
    map[4]=0;
    map[5]=0;
    map[6]=0;
    map[7]=0;
    map[8]=0;
    map[9]=0;
    map[10]=0;
    map[11]=0;
    map[12]=0;
    map[13]=0;
    map[14]=0;
    map[15]=0;
    map[16]=0;
    map[17]=0;
    map[18]=0;
    map[19]=0;
    map[20]=0;
    map[21]=0;
    map[22]=0;
    map[23]=0;
    map[24]=0;
    map[25]=0;
    map[26]=0;
    map[27]=0;
    map[28]=0;
    map[29]=0;
    map[30]=1;
    map[31]=1;
    map[32]=1;
    map[33]=1;
    map[34]=1;
    map[35]=1;
    map[36]=1;
    map[37]=1;
    map[38]=1;
    map[39]=1;
    map[40]=1;
    map[41]=1;
    map[42]=1;
    map[43]=0;
    map[44]=1;
    map[45]=1;
    map[46]=1;
    map[47]=1;
    map[48]=1;
    map[49]=1;
    map[50]=1;
    map[51]=1;
    map[52]=1;
    map[53]=1;
    map[54]=1;
    map[55]=1;
    map[56]=1;
    map[57]=0;
    map[58]=0;
    map[59]=1;
    map[60]=1;
    map[61]=1;
    map[62]=1;
    map[63]=1;
    map[64]=1;
    map[65]=1;
    map[66]=1;
    map[67]=1;
    map[68]=1;
    map[69]=1;
    map[70]=1;
    map[71]=1;
    map[72]=0;
    map[73]=1;
    map[74]=1;
    map[75]=1;
    map[76]=1;
    map[77]=1;
    map[78]=1;
    map[79]=1;
    map[80]=1;
    map[81]=1;
    map[82]=1;
    map[83]=1;
    map[84]=1;
    map[85]=1;
    map[86]=0;
    map[87]=0;
    map[88]=1;
    map[89]=1;
    map[90]=0;
    map[91]=0;
    map[92]=0;
    map[93]=1;
    map[94]=1;
    map[95]=0;
    map[96]=0;
    map[97]=0;
    map[98]=0;
    map[99]=1;
    map[100]=1;
    map[101]=0;
    map[102]=1;
    map[103]=1;
    map[104]=0;
    map[105]=0;
    map[106]=0;
    map[107]=0;
    map[108]=1;
    map[109]=1;
    map[110]=0;
    map[111]=0;
    map[112]=0;
    map[113]=1;
    map[114]=1;
    map[115]=0;
    map[116]=0;
    map[117]=1;
    map[118]=1;
    map[119]=0;
    map[120]=0;
    map[121]=0;
    map[122]=1;
    map[123]=1;
    map[124]=0;
    map[125]=0;
    map[126]=0;
    map[127]=0;
    map[128]=1;
    map[129]=1;
    map[130]=0;
    map[131]=1;
    map[132]=1;
    map[133]=0;
    map[134]=0;
    map[135]=0;
    map[136]=0;
    map[137]=1;
    map[138]=1;
    map[139]=0;
    map[140]=0;
    map[141]=0;
    map[142]=1;
    map[143]=1;
    map[144]=0;
    map[145]=0;
    map[146]=1;
    map[147]=1;
    map[148]=1;
    map[149]=1;
    map[150]=1;
    map[151]=1;
    map[152]=1;
    map[153]=1;
    map[154]=1;
    map[155]=1;
    map[156]=1;
    map[157]=1;
    map[158]=1;
    map[159]=1;
    map[160]=1;
    map[161]=1;
    map[162]=1;
    map[163]=1;
    map[164]=1;
    map[165]=1;
    map[166]=1;
    map[167]=1;
    map[168]=1;
    map[169]=1;
    map[170]=1;
    map[171]=1;
    map[172]=1;
    map[173]=0;
    map[174]=0;
    map[175]=1;
    map[176]=1;
    map[177]=1;
    map[178]=1;
    map[179]=1;
    map[180]=1;
    map[181]=1;
    map[182]=1;
    map[183]=1;
    map[184]=1;
    map[185]=1;
    map[186]=1;
    map[187]=1;
    map[188]=1;
    map[189]=1;
    map[190]=1;
    map[191]=1;
    map[192]=1;
    map[193]=1;
    map[194]=1;
    map[195]=1;
    map[196]=1;
    map[197]=1;
    map[198]=1;
    map[199]=1;
    map[200]=1;
    map[201]=1;
    map[202]=0;
    map[203]=0;
    map[204]=1;
    map[205]=1;
    map[206]=0;
    map[207]=0;
    map[208]=0;
    map[209]=1;
    map[210]=1;
    map[211]=0;
    map[212]=1;
    map[213]=1;
    map[214]=0;
    map[215]=0;
    map[216]=0;
    map[217]=0;
    map[218]=0;
    map[219]=0;
    map[220]=0;
    map[221]=1;
    map[222]=1;
    map[223]=0;
    map[224]=1;
    map[225]=1;
    map[226]=0;
    map[227]=0;
    map[228]=0;
    map[229]=1;
    map[230]=1;
    map[231]=0;
    map[232]=0;
    map[233]=1;
    map[234]=1;
    map[235]=1;
    map[236]=1;
    map[237]=1;
    map[238]=1;
    map[239]=1;
    map[240]=0;
    map[241]=1;
    map[242]=1;
    map[243]=1;
    map[244]=1;
    map[245]=1;
    map[246]=0;
    map[247]=1;
    map[248]=1;
    map[249]=1;
    map[250]=1;
    map[251]=1;
    map[252]=0;
    map[253]=1;
    map[254]=1;
    map[255]=1;
    map[256]=1;
    map[257]=1;
    map[258]=1;
    map[259]=1;
    map[260]=0;
    map[261]=0;
    map[262]=1;
    map[263]=1;
    map[264]=1;
    map[265]=1;
    map[266]=1;
    map[267]=1;
    map[268]=1;
    map[269]=0;
    map[270]=1;
    map[271]=1;
    map[272]=1;
    map[273]=1;
    map[274]=1;
    map[275]=0;
    map[276]=1;
    map[277]=1;
    map[278]=1;
    map[279]=1;
    map[280]=1;
    map[281]=0;
    map[282]=1;
    map[283]=1;
    map[284]=1;
    map[285]=1;
    map[286]=1;
    map[287]=1;
    map[288]=1;
    map[289]=0;
    map[290]=0;
    map[291]=0;
    map[292]=0;
    map[293]=0;
    map[294]=0;
    map[295]=0;
    map[296]=1;
    map[297]=1;
    map[298]=0;
    map[299]=0;
    map[300]=0;
    map[301]=0;
    map[302]=1;
    map[303]=1;
    map[304]=0;
    map[305]=1;
    map[306]=1;
    map[307]=0;
    map[308]=0;
    map[309]=0;
    map[310]=0;
    map[311]=1;
    map[312]=1;
    map[313]=0;
    map[314]=0;
    map[315]=0;
    map[316]=0;
    map[317]=0;
    map[318]=0;
    map[319]=1;
    map[320]=1;
    map[321]=1;
    map[322]=1;
    map[323]=1;
    map[324]=0;
    map[325]=1;
    map[326]=1;
    map[327]=0;
    map[328]=1;
    map[329]=1;
    map[330]=1;
    map[331]=1;
    map[332]=1;
    map[333]=1;
    map[334]=1;
    map[335]=1;
    map[336]=1;
    map[337]=1;
    map[338]=1;
    map[339]=0;
    map[340]=1;
    map[341]=1;
    map[342]=0;
    map[343]=1;
    map[344]=1;
    map[345]=1;
    map[346]=1;
    map[347]=1;
    map[348]=1;
    map[349]=1;
    map[350]=1;
    map[351]=1;
    map[352]=1;
    map[353]=0;
    map[354]=1;
    map[355]=1;
    map[356]=0;
    map[357]=1;
    map[358]=1;
    map[359]=1;
    map[360]=1;
    map[361]=1;
    map[362]=1;
    map[363]=1;
    map[364]=1;
    map[365]=1;
    map[366]=1;
    map[367]=1;
    map[368]=0;
    map[369]=1;
    map[370]=1;
    map[371]=0;
    map[372]=1;
    map[373]=1;
    map[374]=1;
    map[375]=1;
    map[376]=1;
    map[377]=1;
    map[378]=1;
    map[379]=1;
    map[380]=1;
    map[381]=1;
    map[382]=0;
    map[383]=1;
    map[384]=1;
    map[385]=0;
    map[386]=1;
    map[387]=1;
    map[388]=0;
    map[389]=0;
    map[390]=1;
    map[391]=1;
    map[392]=1;
    map[393]=0;
    map[394]=0;
    map[395]=1;
    map[396]=1;
    map[397]=0;
    map[398]=1;
    map[399]=1;
    map[400]=0;
    map[401]=1;
    map[402]=1;
    map[403]=1;
    map[404]=1;
    map[405]=1;
    map[406]=0;
    map[407]=0;
    map[408]=0;
    map[409]=0;
    map[410]=0;
    map[411]=0;
    map[412]=1;
    map[413]=1;
    map[414]=1;
    map[415]=1;
    map[416]=1;
    map[417]=0;
    map[418]=1;
    map[419]=1;
    map[420]=1;
    map[421]=1;
    map[422]=1;
    map[423]=0;
    map[424]=1;
    map[425]=1;
    map[426]=1;
    map[427]=1;
    map[428]=1;
    map[429]=0;
    map[430]=0;
    map[431]=0;
    map[432]=0;
    map[433]=0;
    map[434]=0;
    map[435]=1;
    map[436]=1;
    map[437]=1;
    map[438]=1;
    map[439]=1;
    map[440]=1;
    map[441]=1;
    map[442]=1;
    map[443]=1;
    map[444]=1;
    map[445]=1;
    map[446]=0;
    map[447]=1;
    map[448]=1;
    map[449]=1;
    map[450]=1;
    map[451]=1;
    map[452]=0;
    map[453]=1;
    map[454]=1;
    map[455]=1;
    map[456]=1;
    map[457]=1;
    map[458]=1;
    map[459]=1;
    map[460]=1;
    map[461]=1;
    map[462]=1;
    map[463]=1;
    map[464]=1;
    map[465]=1;
    map[466]=1;
    map[467]=1;
    map[468]=1;
    map[469]=1;
    map[470]=1;
    map[471]=1;
    map[472]=1;
    map[473]=1;
    map[474]=1;
    map[475]=0;
    map[476]=1;
    map[477]=1;
    map[478]=1;
    map[479]=1;
    map[480]=1;
    map[481]=0;
    map[482]=1;
    map[483]=1;
    map[484]=1;
    map[485]=1;
    map[486]=1;
    map[487]=1;
    map[488]=1;
    map[489]=1;
    map[490]=1;
    map[491]=1;
    map[492]=1;
    map[493]=0;
    map[494]=0;
    map[495]=0;
    map[496]=0;
    map[497]=0;
    map[498]=0;
    map[499]=1;
    map[500]=1;
    map[501]=0;
    map[502]=1;
    map[503]=1;
    map[504]=0;
    map[505]=0;
    map[506]=0;
    map[507]=0;
    map[508]=0;
    map[509]=0;
    map[510]=0;
    map[511]=1;
    map[512]=1;
    map[513]=0;
    map[514]=1;
    map[515]=1;
    map[516]=0;
    map[517]=0;
    map[518]=0;
    map[519]=0;
    map[520]=0;
    map[521]=0;
    map[522]=1;
    map[523]=1;
    map[524]=1;
    map[525]=1;
    map[526]=1;
    map[527]=0;
    map[528]=1;
    map[529]=1;
    map[530]=0;
    map[531]=1;
    map[532]=1;
    map[533]=1;
    map[534]=1;
    map[535]=1;
    map[536]=1;
    map[537]=1;
    map[538]=1;
    map[539]=1;
    map[540]=1;
    map[541]=1;
    map[542]=0;
    map[543]=1;
    map[544]=1;
    map[545]=0;
    map[546]=1;
    map[547]=1;
    map[548]=1;
    map[549]=1;
    map[550]=1;
    map[551]=1;
    map[552]=1;
    map[553]=1;
    map[554]=1;
    map[555]=1;
    map[556]=0;
    map[557]=1;
    map[558]=1;
    map[559]=0;
    map[560]=1;
    map[561]=1;
    map[562]=1;
    map[563]=1;
    map[564]=1;
    map[565]=1;
    map[566]=1;
    map[567]=1;
    map[568]=1;
    map[569]=1;
    map[570]=1;
    map[571]=0;
    map[572]=1;
    map[573]=1;
    map[574]=0;
    map[575]=1;
    map[576]=1;
    map[577]=1;
    map[578]=1;
    map[579]=1;
    map[580]=1;
    map[581]=1;
    map[582]=1;
    map[583]=1;
    map[584]=1;
    map[585]=0;
    map[586]=1;
    map[587]=1;
    map[588]=0;
    map[589]=1;
    map[590]=1;
    map[591]=1;
    map[592]=1;
    map[593]=1;
    map[594]=1;
    map[595]=1;
    map[596]=1;
    map[597]=1;
    map[598]=1;
    map[599]=1;
    map[600]=0;
    map[601]=1;
    map[602]=1;
    map[603]=0;
    map[604]=1;
    map[605]=1;
    map[606]=1;
    map[607]=1;
    map[608]=1;
    map[609]=0;
    map[610]=0;
    map[611]=0;
    map[612]=0;
    map[613]=0;
    map[614]=0;
    map[615]=1;
    map[616]=1;
    map[617]=0;
    map[618]=1;
    map[619]=1;
    map[620]=0;
    map[621]=0;
    map[622]=0;
    map[623]=0;
    map[624]=0;
    map[625]=0;
    map[626]=0;
    map[627]=1;
    map[628]=1;
    map[629]=0;
    map[630]=1;
    map[631]=1;
    map[632]=0;
    map[633]=0;
    map[634]=0;
    map[635]=0;
    map[636]=0;
    map[637]=0;
    map[638]=0;
    map[639]=1;
    map[640]=1;
    map[641]=1;
    map[642]=1;
    map[643]=1;
    map[644]=1;
    map[645]=1;
    map[646]=1;
    map[647]=1;
    map[648]=1;
    map[649]=1;
    map[650]=1;
    map[651]=1;
    map[652]=0;
    map[653]=1;
    map[654]=1;
    map[655]=1;
    map[656]=1;
    map[657]=1;
    map[658]=1;
    map[659]=1;
    map[660]=1;
    map[661]=1;
    map[662]=1;
    map[663]=1;
    map[664]=1;
    map[665]=1;
    map[666]=0;
    map[667]=0;
    map[668]=1;
    map[669]=1;
    map[670]=1;
    map[671]=1;
    map[672]=1;
    map[673]=1;
    map[674]=1;
    map[675]=1;
    map[676]=1;
    map[677]=1;
    map[678]=1;
    map[679]=1;
    map[680]=1;
    map[681]=0;
    map[682]=1;
    map[683]=1;
    map[684]=1;
    map[685]=1;
    map[686]=1;
    map[687]=1;
    map[688]=1;
    map[689]=1;
    map[690]=1;
    map[691]=1;
    map[692]=1;
    map[693]=1;
    map[694]=1;
    map[695]=0;
    map[696]=0;
    map[697]=1;
    map[698]=1;
    map[699]=0;
    map[700]=0;
    map[701]=0;
    map[702]=1;
    map[703]=1;
    map[704]=0;
    map[705]=0;
    map[706]=0;
    map[707]=0;
    map[708]=1;
    map[709]=1;
    map[710]=0;
    map[711]=1;
    map[712]=1;
    map[713]=0;
    map[714]=0;
    map[715]=0;
    map[716]=0;
    map[717]=1;
    map[718]=1;
    map[719]=0;
    map[720]=0;
    map[721]=0;
    map[722]=1;
    map[723]=1;
    map[724]=0;
    map[725]=0;
    map[726]=1;
    map[727]=1;
    map[728]=1;
    map[729]=1;
    map[730]=0;
    map[731]=1;
    map[732]=1;
    map[733]=1;
    map[734]=1;
    map[735]=1;
    map[736]=1;
    map[737]=1;
    map[738]=1;
    map[739]=1;
    map[740]=1;
    map[741]=1;
    map[742]=1;
    map[743]=1;
    map[744]=1;
    map[745]=1;
    map[746]=1;
    map[747]=1;
    map[748]=0;
    map[749]=1;
    map[750]=1;
    map[751]=1;
    map[752]=1;
    map[753]=0;
    map[754]=0;
    map[755]=1;
    map[756]=1;
    map[757]=1;
    map[758]=1;
    map[759]=0;
    map[760]=1;
    map[761]=1;
    map[762]=1;
    map[763]=1;
    map[764]=1;
    map[765]=1;
    map[766]=1;
    map[767]=1;
    map[768]=1;
    map[769]=1;
    map[770]=1;
    map[771]=1;
    map[772]=1;
    map[773]=1;
    map[774]=1;
    map[775]=1;
    map[776]=1;
    map[777]=0;
    map[778]=1;
    map[779]=1;
    map[780]=1;
    map[781]=1;
    map[782]=0;
    map[783]=0;
    map[784]=0;
    map[785]=0;
    map[786]=1;
    map[787]=1;
    map[788]=0;
    map[789]=1;
    map[790]=1;
    map[791]=0;
    map[792]=1;
    map[793]=1;
    map[794]=0;
    map[795]=0;
    map[796]=0;
    map[797]=0;
    map[798]=0;
    map[799]=0;
    map[800]=0;
    map[801]=1;
    map[802]=1;
    map[803]=0;
    map[804]=1;
    map[805]=1;
    map[806]=0;
    map[807]=1;
    map[808]=1;
    map[809]=0;
    map[810]=0;
    map[811]=0;
    map[812]=0;
    map[813]=1;
    map[814]=1;
    map[815]=1;
    map[816]=1;
    map[817]=1;
    map[818]=1;
    map[819]=1;
    map[820]=0;
    map[821]=1;
    map[822]=1;
    map[823]=1;
    map[824]=1;
    map[825]=1;
    map[826]=0;
    map[827]=1;
    map[828]=1;
    map[829]=1;
    map[830]=1;
    map[831]=1;
    map[832]=0;
    map[833]=1;
    map[834]=1;
    map[835]=1;
    map[836]=1;
    map[837]=1;
    map[838]=1;
    map[839]=1;
    map[840]=0;
    map[841]=0;
    map[842]=1;
    map[843]=1;
    map[844]=1;
    map[845]=1;
    map[846]=1;
    map[847]=1;
    map[848]=1;
    map[849]=0;
    map[850]=1;
    map[851]=1;
    map[852]=1;
    map[853]=1;
    map[854]=1;
    map[855]=0;
    map[856]=1;
    map[857]=1;
    map[858]=1;
    map[859]=1;
    map[860]=1;
    map[861]=0;
    map[862]=1;
    map[863]=1;
    map[864]=1;
    map[865]=1;
    map[866]=1;
    map[867]=1;
    map[868]=1;
    map[869]=0;
    map[870]=0;
    map[871]=1;
    map[872]=1;
    map[873]=0;
    map[874]=0;
    map[875]=0;
    map[876]=0;
    map[877]=0;
    map[878]=0;
    map[879]=0;
    map[880]=0;
    map[881]=0;
    map[882]=1;
    map[883]=1;
    map[884]=0;
    map[885]=1;
    map[886]=1;
    map[887]=0;
    map[888]=0;
    map[889]=0;
    map[890]=0;
    map[891]=0;
    map[892]=0;
    map[893]=0;
    map[894]=0;
    map[895]=0;
    map[896]=1;
    map[897]=1;
    map[898]=0;
    map[899]=0;
    map[900]=1;
    map[901]=1;
    map[902]=1;
    map[903]=1;
    map[904]=1;
    map[905]=1;
    map[906]=1;
    map[907]=1;
    map[908]=1;
    map[909]=1;
    map[910]=1;
    map[911]=1;
    map[912]=1;
    map[913]=1;
    map[914]=1;
    map[915]=1;
    map[916]=1;
    map[917]=1;
    map[918]=1;
    map[919]=1;
    map[920]=1;
    map[921]=1;
    map[922]=1;
    map[923]=1;
    map[924]=1;
    map[925]=1;
    map[926]=1;
    map[927]=0;
    map[928]=0;
    map[929]=1;
    map[930]=1;
    map[931]=1;
    map[932]=1;
    map[933]=1;
    map[934]=1;
    map[935]=1;
    map[936]=1;
    map[937]=1;
    map[938]=1;
    map[939]=1;
    map[940]=1;
    map[941]=1;
    map[942]=1;
    map[943]=1;
    map[944]=1;
    map[945]=1;
    map[946]=1;
    map[947]=1;
    map[948]=1;
    map[949]=1;
    map[950]=1;
    map[951]=1;
    map[952]=1;
    map[953]=1;
    map[954]=1;
    map[955]=1;
    map[956]=0;
    map[957]=0;
    map[958]=0;
    map[959]=0;
    map[960]=0;
    map[961]=0;
    map[962]=0;
    map[963]=0;
    map[964]=0;
    map[965]=0;
    map[966]=0;
    map[967]=0;
    map[968]=0;
    map[969]=0;
    map[970]=0;
    map[971]=0;
    map[972]=0;
    map[973]=0;
    map[974]=0;
    map[975]=0;
    map[976]=0;
    map[977]=0;
    map[978]=0;
    map[979]=0;
    map[980]=0;
    map[981]=0;
    map[982]=0;
    map[983]=0;
    map[984]=0;
    map[985]=0;
end

assign dot = map[(query_y / 12) * 29 + (query_x / 12)];

always @(posedge clk)
begin
    if (map[(set_y / 12) * 29 + (set_x / 12)] != 0)
    begin
        new <= 1;
        map[(set_y / 12) * 29 + (set_x / 12)] <= 0;
    end
end

endmodule
