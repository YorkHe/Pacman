module monster_ROM(
    clk,
    x,
    y,
    pixel
);

input clk;
input [5:0] x, y;

output reg [2:0] pixel;

localparam MONSTER = {
    24'd111111110000000011111111,
    24'd111111000000000000111111,
    24'd111110000000000000011111,
    24'd111002222000000222200111,
    24'd111022222200002222220111,
    24'd110223333220022333322011,
    24'd100223333220022333322001,
    24'd000223333220022333322000,
    24'd000223333220022333322000,
    24'd000022222200002222220000,
    24'd000002222000000222200000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd000000000000000000000000,
    24'd100000001000000010000001,
    24'd110000011100000111000011,
    24'd111000111110001111100111
};

always @(posedge clk)
begin
    pixel <= MONSTER[y * 24 + x];
end

endmodule
